module test;
  initial begin
    $display("Verilog is alive.");
    $finish;
  end
endmodule
